module multiplier_32bit(P, A, B);
    input [31:0]	A;
    input [31:0]	B;
    output [63:0]	P;

    wire [31:0]	w0,w1,w3,w4,w6,w7,w9,w10,w12,w13,w15,w16,w18,w19,w21,w22,w24,w25,w27,w28,w30,w31,w33,w34,w36,w37,w39,w40,w42,w43,w45,w46,w48,w49,w51,w52,w54,w55,w57,w58,w60,w61,w63,w64,w66,w67,w69,w70,w72,w73,w75,w76,w78,w79,w81,w82,w84,w85,w87,w88,w90,w91;
    wire [32:0]	w2,w5,w8,w11,w14,w17,w20,w23,w26,w29,w32,w35,w38,w41,w44,w47,w50,w53,w56,w59,w62,w65,w68,w71,w74,w77,w80,w83,w86,w89;

and(P[0],A[0],B[0]);
and(w0[0],A[1],B[0]);
and(w0[1],A[2],B[0]);
and(w0[2],A[3],B[0]);
and(w0[3],A[4],B[0]);
and(w0[4],A[5],B[0]);
and(w0[5],A[6],B[0]);
and(w0[6],A[7],B[0]);
and(w0[7],A[8],B[0]);
and(w0[8],A[9],B[0]);
and(w0[9],A[10],B[0]);
and(w0[10],A[11],B[0]);
and(w0[11],A[12],B[0]);
and(w0[12],A[13],B[0]);
and(w0[13],A[14],B[0]);
and(w0[14],A[15],B[0]);
and(w0[15],A[16],B[0]);
and(w0[16],A[17],B[0]);
and(w0[17],A[18],B[0]);
and(w0[18],A[19],B[0]);
and(w0[19],A[20],B[0]);
and(w0[20],A[21],B[0]);
and(w0[21],A[22],B[0]);
and(w0[22],A[23],B[0]);
and(w0[23],A[24],B[0]);
and(w0[24],A[25],B[0]);
and(w0[25],A[26],B[0]);
and(w0[26],A[27],B[0]);
and(w0[27],A[28],B[0]);
and(w0[28],A[29],B[0]);
and(w0[29],A[30],B[0]);
and(w0[30],A[31],B[0]);
and(w0[31],1'b0,1'b0);

and(w1[0],A[0],B[1]);
and(w1[1],A[1],B[1]);
and(w1[2],A[2],B[1]);
and(w1[3],A[3],B[1]);
and(w1[4],A[4],B[1]);
and(w1[5],A[5],B[1]);
and(w1[6],A[6],B[1]);
and(w1[7],A[7],B[1]);
and(w1[8],A[8],B[1]);
and(w1[9],A[9],B[1]);
and(w1[10],A[10],B[1]);
and(w1[11],A[11],B[1]);
and(w1[12],A[12],B[1]);
and(w1[13],A[13],B[1]);
and(w1[14],A[14],B[1]);
and(w1[15],A[15],B[1]);
and(w1[16],A[16],B[1]);
and(w1[17],A[17],B[1]);
and(w1[18],A[18],B[1]);
and(w1[19],A[19],B[1]);
and(w1[20],A[20],B[1]);
and(w1[21],A[21],B[1]);
and(w1[22],A[22],B[1]);
and(w1[23],A[23],B[1]);
and(w1[24],A[24],B[1]);
and(w1[25],A[25],B[1]);
and(w1[26],A[26],B[1]);
and(w1[27],A[27],B[1]);
and(w1[28],A[28],B[1]);
and(w1[29],A[29],B[1]);
and(w1[30],A[30],B[1]);
and(w1[31],A[31],B[1]);

and(w3[0],A[0],B[2]);
and(w3[1],A[1],B[2]);
and(w3[2],A[2],B[2]);
and(w3[3],A[3],B[2]);
and(w3[4],A[4],B[2]);
and(w3[5],A[5],B[2]);
and(w3[6],A[6],B[2]);
and(w3[7],A[7],B[2]);
and(w3[8],A[8],B[2]);
and(w3[9],A[9],B[2]);
and(w3[10],A[10],B[2]);
and(w3[11],A[11],B[2]);
and(w3[12],A[12],B[2]);
and(w3[13],A[13],B[2]);
and(w3[14],A[14],B[2]);
and(w3[15],A[15],B[2]);
and(w3[16],A[16],B[2]);
and(w3[17],A[17],B[2]);
and(w3[18],A[18],B[2]);
and(w3[19],A[19],B[2]);
and(w3[20],A[20],B[2]);
and(w3[21],A[21],B[2]);
and(w3[22],A[22],B[2]);
and(w3[23],A[23],B[2]);
and(w3[24],A[24],B[2]);
and(w3[25],A[25],B[2]);
and(w3[26],A[26],B[2]);
and(w3[27],A[27],B[2]);
and(w3[28],A[28],B[2]);
and(w3[29],A[29],B[2]);
and(w3[30],A[30],B[2]);
and(w3[31],A[31],B[2]);



and(w6[0],A[0],B[3]);
and(w6[1],A[1],B[3]);
and(w6[2],A[2],B[3]);
and(w6[3],A[3],B[3]);
and(w6[4],A[4],B[3]);
and(w6[5],A[5],B[3]);
and(w6[6],A[6],B[3]);
and(w6[7],A[7],B[3]);
and(w6[8],A[8],B[3]);
and(w6[9],A[9],B[3]);
and(w6[10],A[10],B[3]);
and(w6[11],A[11],B[3]);
and(w6[12],A[12],B[3]);
and(w6[13],A[13],B[3]);
and(w6[14],A[14],B[3]);
and(w6[15],A[15],B[3]);
and(w6[16],A[16],B[3]);
and(w6[17],A[17],B[3]);
and(w6[18],A[18],B[3]);
and(w6[19],A[19],B[3]);
and(w6[20],A[20],B[3]);
and(w6[21],A[21],B[3]);
and(w6[22],A[22],B[3]);
and(w6[23],A[23],B[3]);
and(w6[24],A[24],B[3]);
and(w6[25],A[25],B[3]);
and(w6[26],A[26],B[3]);
and(w6[27],A[27],B[3]);
and(w6[28],A[28],B[3]);
and(w6[29],A[29],B[3]);
and(w6[30],A[30],B[3]);
and(w6[31],A[31],B[3]);


and(w9[0],A[0],B[4]);
and(w9[1],A[1],B[4]);
and(w9[2],A[2],B[4]);
and(w9[3],A[3],B[4]);
and(w9[4],A[4],B[4]);
and(w9[5],A[5],B[4]);
and(w9[6],A[6],B[4]);
and(w9[7],A[7],B[4]);
and(w9[8],A[8],B[4]);
and(w9[9],A[9],B[4]);
and(w9[10],A[10],B[4]);
and(w9[11],A[11],B[4]);
and(w9[12],A[12],B[4]);
and(w9[13],A[13],B[4]);
and(w9[14],A[14],B[4]);
and(w9[15],A[15],B[4]);
and(w9[16],A[16],B[4]);
and(w9[17],A[17],B[4]);
and(w9[18],A[18],B[4]);
and(w9[19],A[19],B[4]);
and(w9[20],A[20],B[4]);
and(w9[21],A[21],B[4]);
and(w9[22],A[22],B[4]);
and(w9[23],A[23],B[4]);
and(w9[24],A[24],B[4]);
and(w9[25],A[25],B[4]);
and(w9[26],A[26],B[4]);
and(w9[27],A[27],B[4]);
and(w9[28],A[28],B[4]);
and(w9[29],A[29],B[4]);
and(w9[30],A[30],B[4]);
and(w9[31],A[31],B[4]);

and(w12[0],A[0],B[5]);
and(w12[1],A[1],B[5]);
and(w12[2],A[2],B[5]);
and(w12[3],A[3],B[5]);
and(w12[4],A[4],B[5]);
and(w12[5],A[5],B[5]);
and(w12[6],A[6],B[5]);
and(w12[7],A[7],B[5]);
and(w12[8],A[8],B[5]);
and(w12[9],A[9],B[5]);
and(w12[10],A[10],B[5]);
and(w12[11],A[11],B[5]);
and(w12[12],A[12],B[5]);
and(w12[13],A[13],B[5]);
and(w12[14],A[14],B[5]);
and(w12[15],A[15],B[5]);
and(w12[16],A[16],B[5]);
and(w12[17],A[17],B[5]);
and(w12[18],A[18],B[5]);
and(w12[19],A[19],B[5]);
and(w12[20],A[20],B[5]);
and(w12[21],A[21],B[5]);
and(w12[22],A[22],B[5]);
and(w12[23],A[23],B[5]);
and(w12[24],A[24],B[5]);
and(w12[25],A[25],B[5]);
and(w12[26],A[26],B[5]);
and(w12[27],A[27],B[5]);
and(w12[28],A[28],B[5]);
and(w12[29],A[29],B[5]);
and(w12[30],A[30],B[5]);
and(w12[31],A[31],B[5]);

and(w15[0],A[0],B[6]);
and(w15[1],A[1],B[6]);
and(w15[2],A[2],B[6]);
and(w15[3],A[3],B[6]);
and(w15[4],A[4],B[6]);
and(w15[5],A[5],B[6]);
and(w15[6],A[6],B[6]);
and(w15[7],A[7],B[6]);
and(w15[8],A[8],B[6]);
and(w15[9],A[9],B[6]);
and(w15[10],A[10],B[6]);
and(w15[11],A[11],B[6]);
and(w15[12],A[12],B[6]);
and(w15[13],A[13],B[6]);
and(w15[14],A[14],B[6]);
and(w15[15],A[15],B[6]);
and(w15[16],A[16],B[6]);
and(w15[17],A[17],B[6]);
and(w15[18],A[18],B[6]);
and(w15[19],A[19],B[6]);
and(w15[20],A[20],B[6]);
and(w15[21],A[21],B[6]);
and(w15[22],A[22],B[6]);
and(w15[23],A[23],B[6]);
and(w15[24],A[24],B[6]);
and(w15[25],A[25],B[6]);
and(w15[26],A[26],B[6]);
and(w15[27],A[27],B[6]);
and(w15[28],A[28],B[6]);
and(w15[29],A[29],B[6]);
and(w15[30],A[30],B[6]);
and(w15[31],A[31],B[6]);

and(w18[0],A[0],B[7]);
and(w18[1],A[1],B[7]);
and(w18[2],A[2],B[7]);
and(w18[3],A[3],B[7]);
and(w18[4],A[4],B[7]);
and(w18[5],A[5],B[7]);
and(w18[6],A[6],B[7]);
and(w18[7],A[7],B[7]);
and(w18[8],A[8],B[7]);
and(w18[9],A[9],B[7]);
and(w18[10],A[10],B[7]);
and(w18[11],A[11],B[7]);
and(w18[12],A[12],B[7]);
and(w18[13],A[13],B[7]);
and(w18[14],A[14],B[7]);
and(w18[15],A[15],B[7]);
and(w18[16],A[16],B[7]);
and(w18[17],A[17],B[7]);
and(w18[18],A[18],B[7]);
and(w18[19],A[19],B[7]);
and(w18[20],A[20],B[7]);
and(w18[21],A[21],B[7]);
and(w18[22],A[22],B[7]);
and(w18[23],A[23],B[7]);
and(w18[24],A[24],B[7]);
and(w18[25],A[25],B[7]);
and(w18[26],A[26],B[7]);
and(w18[27],A[27],B[7]);
and(w18[28],A[28],B[7]);
and(w18[29],A[29],B[7]);
and(w18[30],A[30],B[7]);
and(w18[31],A[31],B[7]);

and(w21[0],A[0],B[8]);
and(w21[1],A[1],B[8]);
and(w21[2],A[2],B[8]);
and(w21[3],A[3],B[8]);
and(w21[4],A[4],B[8]);
and(w21[5],A[5],B[8]);
and(w21[6],A[6],B[8]);
and(w21[7],A[7],B[8]);
and(w21[8],A[8],B[8]);
and(w21[9],A[9],B[8]);
and(w21[10],A[10],B[8]);
and(w21[11],A[11],B[8]);
and(w21[12],A[12],B[8]);
and(w21[13],A[13],B[8]);
and(w21[14],A[14],B[8]);
and(w21[15],A[15],B[8]);
and(w21[16],A[16],B[8]);
and(w21[17],A[17],B[8]);
and(w21[18],A[18],B[8]);
and(w21[19],A[19],B[8]);
and(w21[20],A[20],B[8]);
and(w21[21],A[21],B[8]);
and(w21[22],A[22],B[8]);
and(w21[23],A[23],B[8]);
and(w21[24],A[24],B[8]);
and(w21[25],A[25],B[8]);
and(w21[26],A[26],B[8]);
and(w21[27],A[27],B[8]);
and(w21[28],A[28],B[8]);
and(w21[29],A[29],B[8]);
and(w21[30],A[30],B[8]);
and(w21[31],A[31],B[8]);


and(w24[0],A[0],B[9]);
and(w24[1],A[1],B[9]);
and(w24[2],A[2],B[9]);
and(w24[3],A[3],B[9]);
and(w24[4],A[4],B[9]);
and(w24[5],A[5],B[9]);
and(w24[6],A[6],B[9]);
and(w24[7],A[7],B[9]);
and(w24[8],A[8],B[9]);
and(w24[9],A[9],B[9]);
and(w24[10],A[10],B[9]);
and(w24[11],A[11],B[9]);
and(w24[12],A[12],B[9]);
and(w24[13],A[13],B[9]);
and(w24[14],A[14],B[9]);
and(w24[15],A[15],B[9]);
and(w24[16],A[16],B[9]);
and(w24[17],A[17],B[9]);
and(w24[18],A[18],B[9]);
and(w24[19],A[19],B[9]);
and(w24[20],A[20],B[9]);
and(w24[21],A[21],B[9]);
and(w24[22],A[22],B[9]);
and(w24[23],A[23],B[9]);
and(w24[24],A[24],B[9]);
and(w24[25],A[25],B[9]);
and(w24[26],A[26],B[9]);
and(w24[27],A[27],B[9]);
and(w24[28],A[28],B[9]);
and(w24[29],A[29],B[9]);
and(w24[30],A[30],B[9]);
and(w24[31],A[31],B[9]);

and(w27[0],A[0],B[10]);
and(w27[1],A[1],B[10]);
and(w27[2],A[2],B[10]);
and(w27[3],A[3],B[10]);
and(w27[4],A[4],B[10]);
and(w27[5],A[5],B[10]);
and(w27[6],A[6],B[10]);
and(w27[7],A[7],B[10]);
and(w27[8],A[8],B[10]);
and(w27[9],A[9],B[10]);
and(w27[10],A[10],B[10]);
and(w27[11],A[11],B[10]);
and(w27[12],A[12],B[10]);
and(w27[13],A[13],B[10]);
and(w27[14],A[14],B[10]);
and(w27[15],A[15],B[10]);
and(w27[16],A[16],B[10]);
and(w27[17],A[17],B[10]);
and(w27[18],A[18],B[10]);
and(w27[19],A[19],B[10]);
and(w27[20],A[20],B[10]);
and(w27[21],A[21],B[10]);
and(w27[22],A[22],B[10]);
and(w27[23],A[23],B[10]);
and(w27[24],A[24],B[10]);
and(w27[25],A[25],B[10]);
and(w27[26],A[26],B[10]);
and(w27[27],A[27],B[10]);
and(w27[28],A[28],B[10]);
and(w27[29],A[29],B[10]);
and(w27[30],A[30],B[10]);
and(w27[31],A[31],B[10]);


and(w30[0],A[0],B[11]);
and(w30[1],A[1],B[11]);
and(w30[2],A[2],B[11]);
and(w30[3],A[3],B[11]);
and(w30[4],A[4],B[11]);
and(w30[5],A[5],B[11]);
and(w30[6],A[6],B[11]);
and(w30[7],A[7],B[11]);
and(w30[8],A[8],B[11]);
and(w30[9],A[9],B[11]);
and(w30[10],A[10],B[11]);
and(w30[11],A[11],B[11]);
and(w30[12],A[12],B[11]);
and(w30[13],A[13],B[11]);
and(w30[14],A[14],B[11]);
and(w30[15],A[15],B[11]);
and(w30[16],A[16],B[11]);
and(w30[17],A[17],B[11]);
and(w30[18],A[18],B[11]);
and(w30[19],A[19],B[11]);
and(w30[20],A[20],B[11]);
and(w30[21],A[21],B[11]);
and(w30[22],A[22],B[11]);
and(w30[23],A[23],B[11]);
and(w30[24],A[24],B[11]);
and(w30[25],A[25],B[11]);
and(w30[26],A[26],B[11]);
and(w30[27],A[27],B[11]);
and(w30[28],A[28],B[11]);
and(w30[29],A[29],B[11]);
and(w30[30],A[30],B[11]);
and(w30[31],A[31],B[11]);


and(w33[0],A[0],B[12]);
and(w33[1],A[1],B[12]);
and(w33[2],A[2],B[12]);
and(w33[3],A[3],B[12]);
and(w33[4],A[4],B[12]);
and(w33[5],A[5],B[12]);
and(w33[6],A[6],B[12]);
and(w33[7],A[7],B[12]);
and(w33[8],A[8],B[12]);
and(w33[9],A[9],B[12]);
and(w33[10],A[10],B[12]);
and(w33[11],A[11],B[12]);
and(w33[12],A[12],B[12]);
and(w33[13],A[13],B[12]);
and(w33[14],A[14],B[12]);
and(w33[15],A[15],B[12]);
and(w33[16],A[16],B[12]);
and(w33[17],A[17],B[12]);
and(w33[18],A[18],B[12]);
and(w33[19],A[19],B[12]);
and(w33[20],A[20],B[12]);
and(w33[21],A[21],B[12]);
and(w33[22],A[22],B[12]);
and(w33[23],A[23],B[12]);
and(w33[24],A[24],B[12]);
and(w33[25],A[25],B[12]);
and(w33[26],A[26],B[12]);
and(w33[27],A[27],B[12]);
and(w33[28],A[28],B[12]);
and(w33[29],A[29],B[12]);
and(w33[30],A[30],B[12]);
and(w33[31],A[31],B[12]);

and(w36[0],A[0],B[13]);
and(w36[1],A[1],B[13]);
and(w36[2],A[2],B[13]);
and(w36[3],A[3],B[13]);
and(w36[4],A[4],B[13]);
and(w36[5],A[5],B[13]);
and(w36[6],A[6],B[13]);
and(w36[7],A[7],B[13]);
and(w36[8],A[8],B[13]);
and(w36[9],A[9],B[13]);
and(w36[10],A[10],B[13]);
and(w36[11],A[11],B[13]);
and(w36[12],A[12],B[13]);
and(w36[13],A[13],B[13]);
and(w36[14],A[14],B[13]);
and(w36[15],A[15],B[13]);
and(w36[16],A[16],B[13]);
and(w36[17],A[17],B[13]);
and(w36[18],A[18],B[13]);
and(w36[19],A[19],B[13]);
and(w36[20],A[20],B[13]);
and(w36[21],A[21],B[13]);
and(w36[22],A[22],B[13]);
and(w36[23],A[23],B[13]);
and(w36[24],A[24],B[13]);
and(w36[25],A[25],B[13]);
and(w36[26],A[26],B[13]);
and(w36[27],A[27],B[13]);
and(w36[28],A[28],B[13]);
and(w36[29],A[29],B[13]);
and(w36[30],A[30],B[13]);
and(w36[31],A[31],B[13]);


and(w39[0],A[0],B[14]);
and(w39[1],A[1],B[14]);
and(w39[2],A[2],B[14]);
and(w39[3],A[3],B[14]);
and(w39[4],A[4],B[14]);
and(w39[5],A[5],B[14]);
and(w39[6],A[6],B[14]);
and(w39[7],A[7],B[14]);
and(w39[8],A[8],B[14]);
and(w39[9],A[9],B[14]);
and(w39[10],A[10],B[14]);
and(w39[11],A[11],B[14]);
and(w39[12],A[12],B[14]);
and(w39[13],A[13],B[14]);
and(w39[14],A[14],B[14]);
and(w39[15],A[15],B[14]);
and(w39[16],A[16],B[14]);
and(w39[17],A[17],B[14]);
and(w39[18],A[18],B[14]);
and(w39[19],A[19],B[14]);
and(w39[20],A[20],B[14]);
and(w39[21],A[21],B[14]);
and(w39[22],A[22],B[14]);
and(w39[23],A[23],B[14]);
and(w39[24],A[24],B[14]);
and(w39[25],A[25],B[14]);
and(w39[26],A[26],B[14]);
and(w39[27],A[27],B[14]);
and(w39[28],A[28],B[14]);
and(w39[29],A[29],B[14]);
and(w39[30],A[30],B[14]);
and(w39[31],A[31],B[14]);

and(w42[0],A[0],B[15]);
and(w42[1],A[1],B[15]);
and(w42[2],A[2],B[15]);
and(w42[3],A[3],B[15]);
and(w42[4],A[4],B[15]);
and(w42[5],A[5],B[15]);
and(w42[6],A[6],B[15]);
and(w42[7],A[7],B[15]);
and(w42[8],A[8],B[15]);
and(w42[9],A[9],B[15]);
and(w42[10],A[10],B[15]);
and(w42[11],A[11],B[15]);
and(w42[12],A[12],B[15]);
and(w42[13],A[13],B[15]);
and(w42[14],A[14],B[15]);
and(w42[15],A[15],B[15]);
and(w42[16],A[16],B[15]);
and(w42[17],A[17],B[15]);
and(w42[18],A[18],B[15]);
and(w42[19],A[19],B[15]);
and(w42[20],A[20],B[15]);
and(w42[21],A[21],B[15]);
and(w42[22],A[22],B[15]);
and(w42[23],A[23],B[15]);
and(w42[24],A[24],B[15]);
and(w42[25],A[25],B[15]);
and(w42[26],A[26],B[15]);
and(w42[27],A[27],B[15]);
and(w42[28],A[28],B[15]);
and(w42[29],A[29],B[15]);
and(w42[30],A[30],B[15]);
and(w42[31],A[31],B[15]);

and(w45[0],A[0],B[16]);
and(w45[1],A[1],B[16]);
and(w45[2],A[2],B[16]);
and(w45[3],A[3],B[16]);
and(w45[4],A[4],B[16]);
and(w45[5],A[5],B[16]);
and(w45[6],A[6],B[16]);
and(w45[7],A[7],B[16]);
and(w45[8],A[8],B[16]);
and(w45[9],A[9],B[16]);
and(w45[10],A[10],B[16]);
and(w45[11],A[11],B[16]);
and(w45[12],A[12],B[16]);
and(w45[13],A[13],B[16]);
and(w45[14],A[14],B[16]);
and(w45[15],A[15],B[16]);
and(w45[16],A[16],B[16]);
and(w45[17],A[17],B[16]);
and(w45[18],A[18],B[16]);
and(w45[19],A[19],B[16]);
and(w45[20],A[20],B[16]);
and(w45[21],A[21],B[16]);
and(w45[22],A[22],B[16]);
and(w45[23],A[23],B[16]);
and(w45[24],A[24],B[16]);
and(w45[25],A[25],B[16]);
and(w45[26],A[26],B[16]);
and(w45[27],A[27],B[16]);
and(w45[28],A[28],B[16]);
and(w45[29],A[29],B[16]);
and(w45[30],A[30],B[16]);
and(w45[31],A[31],B[16]);

and(w48[0],A[0],B[17]);
and(w48[1],A[1],B[17]);
and(w48[2],A[2],B[17]);
and(w48[3],A[3],B[17]);
and(w48[4],A[4],B[17]);
and(w48[5],A[5],B[17]);
and(w48[6],A[6],B[17]);
and(w48[7],A[7],B[17]);
and(w48[8],A[8],B[17]);
and(w48[9],A[9],B[17]);
and(w48[10],A[10],B[17]);
and(w48[11],A[11],B[17]);
and(w48[12],A[12],B[17]);
and(w48[13],A[13],B[17]);
and(w48[14],A[14],B[17]);
and(w48[15],A[15],B[17]);
and(w48[16],A[16],B[17]);
and(w48[17],A[17],B[17]);
and(w48[18],A[18],B[17]);
and(w48[19],A[19],B[17]);
and(w48[20],A[20],B[17]);
and(w48[21],A[21],B[17]);
and(w48[22],A[22],B[17]);
and(w48[23],A[23],B[17]);
and(w48[24],A[24],B[17]);
and(w48[25],A[25],B[17]);
and(w48[26],A[26],B[17]);
and(w48[27],A[27],B[17]);
and(w48[28],A[28],B[17]);
and(w48[29],A[29],B[17]);
and(w48[30],A[30],B[17]);
and(w48[31],A[31],B[17]);



and(w51[0],A[0],B[18]);
and(w51[1],A[1],B[18]);
and(w51[2],A[2],B[18]);
and(w51[3],A[3],B[18]);
and(w51[4],A[4],B[18]);
and(w51[5],A[5],B[18]);
and(w51[6],A[6],B[18]);
and(w51[7],A[7],B[18]);
and(w51[8],A[8],B[18]);
and(w51[9],A[9],B[18]);
and(w51[10],A[10],B[18]);
and(w51[11],A[11],B[18]);
and(w51[12],A[12],B[18]);
and(w51[13],A[13],B[18]);
and(w51[14],A[14],B[18]);
and(w51[15],A[15],B[18]);
and(w51[16],A[16],B[18]);
and(w51[17],A[17],B[18]);
and(w51[18],A[18],B[18]);
and(w51[19],A[19],B[18]);
and(w51[20],A[20],B[18]);
and(w51[21],A[21],B[18]);
and(w51[22],A[22],B[18]);
and(w51[23],A[23],B[18]);
and(w51[24],A[24],B[18]);
and(w51[25],A[25],B[18]);
and(w51[26],A[26],B[18]);
and(w51[27],A[27],B[18]);
and(w51[28],A[28],B[18]);
and(w51[29],A[29],B[18]);
and(w51[30],A[30],B[18]);
and(w51[31],A[31],B[18]);


and(w54[0],A[0],B[19]);
and(w54[1],A[1],B[19]);
and(w54[2],A[2],B[19]);
and(w54[3],A[3],B[19]);
and(w54[4],A[4],B[19]);
and(w54[5],A[5],B[19]);
and(w54[6],A[6],B[19]);
and(w54[7],A[7],B[19]);
and(w54[8],A[8],B[19]);
and(w54[9],A[9],B[19]);
and(w54[10],A[10],B[19]);
and(w54[11],A[11],B[19]);
and(w54[12],A[12],B[19]);
and(w54[13],A[13],B[19]);
and(w54[14],A[14],B[19]);
and(w54[15],A[15],B[19]);
and(w54[16],A[16],B[19]);
and(w54[17],A[17],B[19]);
and(w54[18],A[18],B[19]);
and(w54[19],A[19],B[19]);
and(w54[20],A[20],B[19]);
and(w54[21],A[21],B[19]);
and(w54[22],A[22],B[19]);
and(w54[23],A[23],B[19]);
and(w54[24],A[24],B[19]);
and(w54[25],A[25],B[19]);
and(w54[26],A[26],B[19]);
and(w54[27],A[27],B[19]);
and(w54[28],A[28],B[19]);
and(w54[29],A[29],B[19]);
and(w54[30],A[30],B[19]);
and(w54[31],A[31],B[19]);

and(w57[0],A[0],B[20]);
and(w57[1],A[1],B[20]);
and(w57[2],A[2],B[20]);
and(w57[3],A[3],B[20]);
and(w57[4],A[4],B[20]);
and(w57[5],A[5],B[20]);
and(w57[6],A[6],B[20]);
and(w57[7],A[7],B[20]);
and(w57[8],A[8],B[20]);
and(w57[9],A[9],B[20]);
and(w57[10],A[10],B[20]);
and(w57[11],A[11],B[20]);
and(w57[12],A[12],B[20]);
and(w57[13],A[13],B[20]);
and(w57[14],A[14],B[20]);
and(w57[15],A[15],B[20]);
and(w57[16],A[16],B[20]);
and(w57[17],A[17],B[20]);
and(w57[18],A[18],B[20]);
and(w57[19],A[19],B[20]);
and(w57[20],A[20],B[20]);
and(w57[21],A[21],B[20]);
and(w57[22],A[22],B[20]);
and(w57[23],A[23],B[20]);
and(w57[24],A[24],B[20]);
and(w57[25],A[25],B[20]);
and(w57[26],A[26],B[20]);
and(w57[27],A[27],B[20]);
and(w57[28],A[28],B[20]);
and(w57[29],A[29],B[20]);
and(w57[30],A[30],B[20]);
and(w57[31],A[31],B[20]);

and(w60[0],A[0],B[21]);
and(w60[1],A[1],B[21]);
and(w60[2],A[2],B[21]);
and(w60[3],A[3],B[21]);
and(w60[4],A[4],B[21]);
and(w60[5],A[5],B[21]);
and(w60[6],A[6],B[21]);
and(w60[7],A[7],B[21]);
and(w60[8],A[8],B[21]);
and(w60[9],A[9],B[21]);
and(w60[10],A[10],B[21]);
and(w60[11],A[11],B[21]);
and(w60[12],A[12],B[21]);
and(w60[13],A[13],B[21]);
and(w60[14],A[14],B[21]);
and(w60[15],A[15],B[21]);
and(w60[16],A[16],B[21]);
and(w60[17],A[17],B[21]);
and(w60[18],A[18],B[21]);
and(w60[19],A[19],B[21]);
and(w60[20],A[20],B[21]);
and(w60[21],A[21],B[21]);
and(w60[22],A[22],B[21]);
and(w60[23],A[23],B[21]);
and(w60[24],A[24],B[21]);
and(w60[25],A[25],B[21]);
and(w60[26],A[26],B[21]);
and(w60[27],A[27],B[21]);
and(w60[28],A[28],B[21]);
and(w60[29],A[29],B[21]);
and(w60[30],A[30],B[21]);
and(w60[31],A[31],B[21]);

and(w63[0],A[0],B[22]);
and(w63[1],A[1],B[22]);
and(w63[2],A[2],B[22]);
and(w63[3],A[3],B[22]);
and(w63[4],A[4],B[22]);
and(w63[5],A[5],B[22]);
and(w63[6],A[6],B[22]);
and(w63[7],A[7],B[22]);
and(w63[8],A[8],B[22]);
and(w63[9],A[9],B[22]);
and(w63[10],A[10],B[22]);
and(w63[11],A[11],B[22]);
and(w63[12],A[12],B[22]);
and(w63[13],A[13],B[22]);
and(w63[14],A[14],B[22]);
and(w63[15],A[15],B[22]);
and(w63[16],A[16],B[22]);
and(w63[17],A[17],B[22]);
and(w63[18],A[18],B[22]);
and(w63[19],A[19],B[22]);
and(w63[20],A[20],B[22]);
and(w63[21],A[21],B[22]);
and(w63[22],A[22],B[22]);
and(w63[23],A[23],B[22]);
and(w63[24],A[24],B[22]);
and(w63[25],A[25],B[22]);
and(w63[26],A[26],B[22]);
and(w63[27],A[27],B[22]);
and(w63[28],A[28],B[22]);
and(w63[29],A[29],B[22]);
and(w63[30],A[30],B[22]);
and(w63[31],A[31],B[22]);

and(w66[0],A[0],B[23]);
and(w66[1],A[1],B[23]);
and(w66[2],A[2],B[23]);
and(w66[3],A[3],B[23]);
and(w66[4],A[4],B[23]);
and(w66[5],A[5],B[23]);
and(w66[6],A[6],B[23]);
and(w66[7],A[7],B[23]);
and(w66[8],A[8],B[23]);
and(w66[9],A[9],B[23]);
and(w66[10],A[10],B[23]);
and(w66[11],A[11],B[23]);
and(w66[12],A[12],B[23]);
and(w66[13],A[13],B[23]);
and(w66[14],A[14],B[23]);
and(w66[15],A[15],B[23]);
and(w66[16],A[16],B[23]);
and(w66[17],A[17],B[23]);
and(w66[18],A[18],B[23]);
and(w66[19],A[19],B[23]);
and(w66[20],A[20],B[23]);
and(w66[21],A[21],B[23]);
and(w66[22],A[22],B[23]);
and(w66[23],A[23],B[23]);
and(w66[24],A[24],B[23]);
and(w66[25],A[25],B[23]);
and(w66[26],A[26],B[23]);
and(w66[27],A[27],B[23]);
and(w66[28],A[28],B[23]);
and(w66[29],A[29],B[23]);
and(w66[30],A[30],B[23]);
and(w66[31],A[31],B[23]);


and(w69[0],A[0],B[24]);
and(w69[1],A[1],B[24]);
and(w69[2],A[2],B[24]);
and(w69[3],A[3],B[24]);
and(w69[4],A[4],B[24]);
and(w69[5],A[5],B[24]);
and(w69[6],A[6],B[24]);
and(w69[7],A[7],B[24]);
and(w69[8],A[8],B[24]);
and(w69[9],A[9],B[24]);
and(w69[10],A[10],B[24]);
and(w69[11],A[11],B[24]);
and(w69[12],A[12],B[24]);
and(w69[13],A[13],B[24]);
and(w69[14],A[14],B[24]);
and(w69[15],A[15],B[24]);
and(w69[16],A[16],B[24]);
and(w69[17],A[17],B[24]);
and(w69[18],A[18],B[24]);
and(w69[19],A[19],B[24]);
and(w69[20],A[20],B[24]);
and(w69[21],A[21],B[24]);
and(w69[22],A[22],B[24]);
and(w69[23],A[23],B[24]);
and(w69[24],A[24],B[24]);
and(w69[25],A[25],B[24]);
and(w69[26],A[26],B[24]);
and(w69[27],A[27],B[24]);
and(w69[28],A[28],B[24]);
and(w69[29],A[29],B[24]);
and(w69[30],A[30],B[24]);
and(w69[31],A[31],B[24]);

and(w72[0],A[0],B[25]);
and(w72[1],A[1],B[25]);
and(w72[2],A[2],B[25]);
and(w72[3],A[3],B[25]);
and(w72[4],A[4],B[25]);
and(w72[5],A[5],B[25]);
and(w72[6],A[6],B[25]);
and(w72[7],A[7],B[25]);
and(w72[8],A[8],B[25]);
and(w72[9],A[9],B[25]);
and(w72[10],A[10],B[25]);
and(w72[11],A[11],B[25]);
and(w72[12],A[12],B[25]);
and(w72[13],A[13],B[25]);
and(w72[14],A[14],B[25]);
and(w72[15],A[15],B[25]);
and(w72[16],A[16],B[25]);
and(w72[17],A[17],B[25]);
and(w72[18],A[18],B[25]);
and(w72[19],A[19],B[25]);
and(w72[20],A[20],B[25]);
and(w72[21],A[21],B[25]);
and(w72[22],A[22],B[25]);
and(w72[23],A[23],B[25]);
and(w72[24],A[24],B[25]);
and(w72[25],A[25],B[25]);
and(w72[26],A[26],B[25]);
and(w72[27],A[27],B[25]);
and(w72[28],A[28],B[25]);
and(w72[29],A[29],B[25]);
and(w72[30],A[30],B[25]);
and(w72[31],A[31],B[25]);


and(w75[0],A[0],B[26]);
and(w75[1],A[1],B[26]);
and(w75[2],A[2],B[26]);
and(w75[3],A[3],B[26]);
and(w75[4],A[4],B[26]);
and(w75[5],A[5],B[26]);
and(w75[6],A[6],B[26]);
and(w75[7],A[7],B[26]);
and(w75[8],A[8],B[26]);
and(w75[9],A[9],B[26]);
and(w75[10],A[10],B[26]);
and(w75[11],A[11],B[26]);
and(w75[12],A[12],B[26]);
and(w75[13],A[13],B[26]);
and(w75[14],A[14],B[26]);
and(w75[15],A[15],B[26]);
and(w75[16],A[16],B[26]);
and(w75[17],A[17],B[26]);
and(w75[18],A[18],B[26]);
and(w75[19],A[19],B[26]);
and(w75[20],A[20],B[26]);
and(w75[21],A[21],B[26]);
and(w75[22],A[22],B[26]);
and(w75[23],A[23],B[26]);
and(w75[24],A[24],B[26]);
and(w75[25],A[25],B[26]);
and(w75[26],A[26],B[26]);
and(w75[27],A[27],B[26]);
and(w75[28],A[28],B[26]);
and(w75[29],A[29],B[26]);
and(w75[30],A[30],B[26]);
and(w75[31],A[31],B[26]);


and(w78[0],A[0],B[27]);
and(w78[1],A[1],B[27]);
and(w78[2],A[2],B[27]);
and(w78[3],A[3],B[27]);
and(w78[4],A[4],B[27]);
and(w78[5],A[5],B[27]);
and(w78[6],A[6],B[27]);
and(w78[7],A[7],B[27]);
and(w78[8],A[8],B[27]);
and(w78[9],A[9],B[27]);
and(w78[10],A[10],B[27]);
and(w78[11],A[11],B[27]);
and(w78[12],A[12],B[27]);
and(w78[13],A[13],B[27]);
and(w78[14],A[14],B[27]);
and(w78[15],A[15],B[27]);
and(w78[16],A[16],B[27]);
and(w78[17],A[17],B[27]);
and(w78[18],A[18],B[27]);
and(w78[19],A[19],B[27]);
and(w78[20],A[20],B[27]);
and(w78[21],A[21],B[27]);
and(w78[22],A[22],B[27]);
and(w78[23],A[23],B[27]);
and(w78[24],A[24],B[27]);
and(w78[25],A[25],B[27]);
and(w78[26],A[26],B[27]);
and(w78[27],A[27],B[27]);
and(w78[28],A[28],B[27]);
and(w78[29],A[29],B[27]);
and(w78[30],A[30],B[27]);
and(w78[31],A[31],B[27]);

and(w81[0],A[0],B[28]);
and(w81[1],A[1],B[28]);
and(w81[2],A[2],B[28]);
and(w81[3],A[3],B[28]);
and(w81[4],A[4],B[28]);
and(w81[5],A[5],B[28]);
and(w81[6],A[6],B[28]);
and(w81[7],A[7],B[28]);
and(w81[8],A[8],B[28]);
and(w81[9],A[9],B[28]);
and(w81[10],A[10],B[28]);
and(w81[11],A[11],B[28]);
and(w81[12],A[12],B[28]);
and(w81[13],A[13],B[28]);
and(w81[14],A[14],B[28]);
and(w81[15],A[15],B[28]);
and(w81[16],A[16],B[28]);
and(w81[17],A[17],B[28]);
and(w81[18],A[18],B[28]);
and(w81[19],A[19],B[28]);
and(w81[20],A[20],B[28]);
and(w81[21],A[21],B[28]);
and(w81[22],A[22],B[28]);
and(w81[23],A[23],B[28]);
and(w81[24],A[24],B[28]);
and(w81[25],A[25],B[28]);
and(w81[26],A[26],B[28]);
and(w81[27],A[27],B[28]);
and(w81[28],A[28],B[28]);
and(w81[29],A[29],B[28]);
and(w81[30],A[30],B[28]);
and(w81[31],A[31],B[28]);


and(w84[0],A[0],B[29]);
and(w84[1],A[1],B[29]);
and(w84[2],A[2],B[29]);
and(w84[3],A[3],B[29]);
and(w84[4],A[4],B[29]);
and(w84[5],A[5],B[29]);
and(w84[6],A[6],B[29]);
and(w84[7],A[7],B[29]);
and(w84[8],A[8],B[29]);
and(w84[9],A[9],B[29]);
and(w84[10],A[10],B[29]);
and(w84[11],A[11],B[29]);
and(w84[12],A[12],B[29]);
and(w84[13],A[13],B[29]);
and(w84[14],A[14],B[29]);
and(w84[15],A[15],B[29]);
and(w84[16],A[16],B[29]);
and(w84[17],A[17],B[29]);
and(w84[18],A[18],B[29]);
and(w84[19],A[19],B[29]);
and(w84[20],A[20],B[29]);
and(w84[21],A[21],B[29]);
and(w84[22],A[22],B[29]);
and(w84[23],A[23],B[29]);
and(w84[24],A[24],B[29]);
and(w84[25],A[25],B[29]);
and(w84[26],A[26],B[29]);
and(w84[27],A[27],B[29]);
and(w84[28],A[28],B[29]);
and(w84[29],A[29],B[29]);
and(w84[30],A[30],B[29]);
and(w84[31],A[31],B[29]);

and(w87[0],A[0],B[30]);
and(w87[1],A[1],B[30]);
and(w87[2],A[2],B[30]);
and(w87[3],A[3],B[30]);
and(w87[4],A[4],B[30]);
and(w87[5],A[5],B[30]);
and(w87[6],A[6],B[30]);
and(w87[7],A[7],B[30]);
and(w87[8],A[8],B[30]);
and(w87[9],A[9],B[30]);
and(w87[10],A[10],B[30]);
and(w87[11],A[11],B[30]);
and(w87[12],A[12],B[30]);
and(w87[13],A[13],B[30]);
and(w87[14],A[14],B[30]);
and(w87[15],A[15],B[30]);
and(w87[16],A[16],B[30]);
and(w87[17],A[17],B[30]);
and(w87[18],A[18],B[30]);
and(w87[19],A[19],B[30]);
and(w87[20],A[20],B[30]);
and(w87[21],A[21],B[30]);
and(w87[22],A[22],B[30]);
and(w87[23],A[23],B[30]);
and(w87[24],A[24],B[30]);
and(w87[25],A[25],B[30]);
and(w87[26],A[26],B[30]);
and(w87[27],A[27],B[30]);
and(w87[28],A[28],B[30]);
and(w87[29],A[29],B[30]);
and(w87[30],A[30],B[30]);
and(w87[31],A[31],B[30]);

and(w90[0],A[0],B[31]);
and(w90[1],A[1],B[31]);
and(w90[2],A[2],B[31]);
and(w90[3],A[3],B[31]);
and(w90[4],A[4],B[31]);
and(w90[5],A[5],B[31]);
and(w90[6],A[6],B[31]);
and(w90[7],A[7],B[31]);
and(w90[8],A[8],B[31]);
and(w90[9],A[9],B[31]);
and(w90[10],A[10],B[31]);
and(w90[11],A[11],B[31]);
and(w90[12],A[12],B[31]);
and(w90[13],A[13],B[31]);
and(w90[14],A[14],B[31]);
and(w90[15],A[15],B[31]);
and(w90[16],A[16],B[31]);
and(w90[17],A[17],B[31]);
and(w90[18],A[18],B[31]);
and(w90[19],A[19],B[31]);
and(w90[20],A[20],B[31]);
and(w90[21],A[21],B[31]);
and(w90[22],A[22],B[31]);
and(w90[23],A[23],B[31]);
and(w90[24],A[24],B[31]);
and(w90[25],A[25],B[31]);
and(w90[26],A[26],B[31]);
and(w90[27],A[27],B[31]);
and(w90[28],A[28],B[31]);
and(w90[29],A[29],B[31]);
and(w90[30],A[30],B[31]);
and(w90[31],A[31],B[31]);


assign P[1]= w2[0];
assign w4[30:0]=w2[31:1];
assign w4[31]=w2[32];

assign P[2]= w5[0];
assign w7[30:0]=w5[31:1];
assign w7[31]=w5[32];

assign P[3]= w8[0];
assign w10[30:0]=w8[31:1];
assign w10[31]=w8[32];

assign P[4]= w11[0];
assign w13[30:0]=w11[31:1];
assign w13[31]=w11[32];

assign P[5]= w14[0];
assign w16[30:0]=w14[31:1];
assign w16[31]=w14[32];

assign P[6]= w17[0];
assign w19[30:0]=w17[31:1];
assign w19[31]=w17[32];

assign P[7]= w20[0];
assign w22[30:0]=w20[31:1];
assign w22[31]=w20[32];

assign P[8]= w23[0];
assign w25[30:0]=w23[31:1];
assign w25[31]=w23[32];

assign P[9]= w26[0];
assign w28[30:0]=w26[31:1];
assign w28[31]=w26[32];

assign P[10]= w29[0];
assign w31[30:0]=w29[31:1];
assign w31[31]=w29[32];

assign P[11]= w32[0];
assign w34[30:0]=w32[31:1];
assign w34[31]=w32[32];

assign P[12]= w35[0];
assign w37[30:0]=w35[31:1];
assign w37[31]=w35[32];

assign P[13]= w38[0];
assign w40[30:0]=w38[31:1];
assign w40[31]=w38[32];

assign P[14]= w41[0];
assign w43[30:0]=w41[31:1];
assign w43[31]=w41[32];

assign P[15]= w44[0];
assign w46[30:0]=w44[31:1];
assign w46[31]=w44[32];

assign P[16]= w47[0];
assign w49[30:0]=w47[31:1];
assign w49[31]=w47[32];

assign P[17]= w50[0];
assign w52[30:0]=w50[31:1];
assign w52[31]=w50[32];

assign P[18]= w53[0];
assign w55[30:0]=w53[31:1];
assign w55[31]=w53[32];

assign P[19]= w56[0];
assign w58[30:0]=w56[31:1];
assign w58[31]=w56[32];

assign P[20]= w59[0];
assign w61[30:0]=w59[31:1];
assign w61[31]=w59[32];

assign P[21]= w62[0];
assign w64[30:0]=w62[31:1];
assign w64[31]=w62[32];

assign P[22]= w65[0];
assign w67[30:0]=w65[31:1];
assign w67[31]=w65[32];

assign P[23]= w68[0];
assign w70[30:0]=w68[31:1];
assign w70[31]=w68[32];

assign P[24]= w71[0];
assign w73[30:0]=w71[31:1];
assign w73[31]=w71[32];

assign P[25]= w74[0];
assign w76[30:0]=w74[31:1];
assign w76[31]=w74[32];

assign P[26]= w77[0];
assign w79[30:0]=w77[31:1];
assign w79[31]=w77[32];

assign P[27]= w80[0];
assign w82[30:0]=w80[31:1];
assign w82[31]=w80[32];

assign P[28]= w83[0];
assign w85[30:0]=w83[31:1];
assign w85[31]=w83[32];

assign P[29]= w86[0];
assign w88[30:0]=w86[31:1];
assign w88[31]=w86[32];

assign P[30]= w89[0];
assign w91[30:0]=w89[31:1];
assign w91[31]=w89[32];

adder_32bit add1(w2[32],w2[31:0],w1,w0,0);
adder_32bit add2(w5[32],w5[31:0],w4,w3,0);
adder_32bit add3(w8[32],w8[31:0],w7,w6,0);
adder_32bit add4(w11[32],w11[31:0],w10,w9,0);
adder_32bit add5(w14[32],w14[31:0],w13,w12,0);
adder_32bit add6(w17[32],w17[31:0],w16,w15,0);
adder_32bit add7(w20[32],w20[31:0],w19,w18,0);
adder_32bit add8(w23[32],w23[31:0],w22,w21,0);
adder_32bit add9(w26[32],w26[31:0],w25,w24,0);
adder_32bit add10(w29[32],w29[31:0],w28,w27,0);
adder_32bit add11(w32[32],w32[31:0],w31,w30,0);
adder_32bit add12(w35[32],w35[31:0],w34,w33,0);
adder_32bit add13(w38[32],w38[31:0],w37,w36,0);
adder_32bit add14(w41[32],w41[31:0],w40,w39,0);
adder_32bit add15(w44[32],w44[31:0],w43,w42,0);
adder_32bit add16(w47[32],w47[31:0],w46,w45,0);
adder_32bit add17(w50[32],w50[31:0],w49,w48,0);
adder_32bit add18(w53[32],w53[31:0],w52,w51,0);
adder_32bit add19(w56[32],w56[31:0],w55,w54,0);
adder_32bit add20(w59[32],w59[31:0],w58,w57,0);
adder_32bit add21(w62[32],w62[31:0],w61,w60,0);
adder_32bit add22(w65[32],w65[31:0],w64,w63,0);
adder_32bit add23(w68[32],w68[31:0],w67,w66,0);
adder_32bit add24(w71[32],w71[31:0],w70,w69,0);
adder_32bit add25(w74[32],w74[31:0],w73,w72,0);
adder_32bit add26(w77[32],w77[31:0],w76,w75,0);
adder_32bit add27(w80[32],w80[31:0],w79,w78,0);
adder_32bit add28(w83[32],w83[31:0],w82,w81,0);
adder_32bit add29(w86[32],w86[31:0],w85,w84,0);
adder_32bit add30(w89[32],w89[31:0],w88,w87,0);
adder_32bit add31(P[63],P[62:31],w91,w90,0);



endmodule
